Diode Characteristic

v1 1 0 0
d1 1 0 dio1
.model dio1 d
.dc v1 0 0.9 0.01  ; ONLY WORKS AFTER run !!! 

.control
* dc v1 0 0.9 0.01
* plot -i(v1)
run
plot -i(v1)
.endc
.end