Basic RC circuit
r 1 2 1.0
c 2 3 1.0u
l 3 0 1.0u
$$$$ l 2 0 1.0e-3
vin 1 0 dc 0 ac 1   $ < the ac source
$$$$ vin 1 0 0.001 ac sin(0  1  1meg)
.options noacct
.ac dec 10 .01 1e6
$$$$ .tran 1ns 5us
.plot ac vdb(2) xlog
.print mag(v(2))
.end
