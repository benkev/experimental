*
* Test IRFD9120 characteristics
*
 
.model IRFD9120 PMOS (Level=3 Gamma=0 Delta=0 Eta=0 Theta=0 Kappa=0.2 Vmax=0 Xj=0 Tox=100n Uo=300 Phi=.6 Rs=.1474 Kp=10.35u W=.29 L=2u Vto=-3.386 Rd=.2494 Rds=444.4K Cbd=899.2p Pb=.8 Mj=.5 Fc=.5 Cgso=5.218n Cgdo=324.8p Rg=7.061 Is=2.618E-18 N=2 Tt=320n)

M1 0 2 1 1 IRFD9120

VDS 1 0 10V
VGS 2 0 2.8V

.dc   VDS  0.001  20  0.1     VGS  6   0.2


.control
set color0=white
run

plot  -i(VDS)
plot loglog -i(VDS)
.endc