Test the BFT46 JFET
* Power
Vdd  2  0  DC  4.0V
* Circuit description
J1  2  1  1  BFT46  ; Jxxx D G S model_name
R1  1  0  100
.MODEL  BFT46   NJF
+             VTO = -6.4188E-001
* +            BETA = 1.86172E-003
+            BETA = 0.5E-003
+          LAMBDA = 2.16604E-002
+              RD = 9.23044E+000
+              RS = 9.23044E+000
+              IS = 1.68833E-016
+            CGS  = 2.20000E-012
+            CGD  = 2.20000E-012
+              PB = 8.27713E-001
+              FC = 5.00000E-001

* .tran  10us  5ms  ; time_step time_stop
.dc Vdd  0  5  0.1
