RC Circuit Transient Responce

r1 1 2 1k
c1 2 0 1u

* pwl: t=0 0V; t=10ms, 0V; t=11ms, 5V; t=20ms, 5V:
vin 1 0 pwl (0 0 10ms 0 11ms 5v); Piecewise Linear

* Transient analysis: step  0.02ms, maximum 20ms
* .tran 0.02ms 20ms

.dc vin  0  5  0.1

.control
run
* plot v(1) v(2)
plot v(2)
set color0=white
set color1=black
set color2=blue
set color3=red
set xbrushwidth=2
* print v(2)
* print v(2) > v_2.txt
* plot v(2) - v(1)
.endc

.end

