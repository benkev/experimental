Compression effect in a JFET amplifier circuit
* Power
Vdd  3  0  DC  4.0V
* Input waveform generator
Vin  1  0  sin(0V  50mV  1000Hz)
* Circuit description
J1  3  2  2  BFT46  ; Jxxx D G S model_name
J2  2  1  0  BFT46  ; Jxxx D G S model_name
R1  1  0  470k
* .model BFT46  NJF  (beta=0.14m Vto=-1.2V lambda=1e-3 Rd=100 Rs=100)
*PHILIPS SEMICONDUCTORS        Version: 1.0
*Filename: BFT46.PRM         Date: Oct 1992
.MODEL  BFT46   NJF
+             VTO = -6.4188E-001
* +            BETA = 1.86172E-003
+            BETA = 0.5E-003
+          LAMBDA = 2.16604E-002
+              RD = 9.23044E+000
+              RS = 9.23044E+000
+              IS = 1.68833E-016
+            CGS  = 2.20000E-012
+            CGD  = 2.20000E-012
+              PB = 8.27713E-001
+              FC = 5.00000E-001

.tran  10us  5ms  ; time_step time_stop

